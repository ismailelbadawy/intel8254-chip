`include "read-write.v"
module rw_tb();

    // we need to test this.
    
endmodule