module counter(input clk, input gate, output reg out);
    // Insert code here.
    
endmodule