module CWR ();


endmodule