module counter()
    // Insert code here.
endmodule